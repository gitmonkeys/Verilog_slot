module finaldesign { input reset, clk, lever,
                     output [7:0] Anode_Activate,
                     output [
