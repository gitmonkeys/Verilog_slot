module clock_divider { input clk, reset,
                       output reg sclk
                     };
  
